`include "common.sv"
`include "inter.sv"
`include "mem.sv"
`include "mem_tx.sv"
`include "gen.sv"
`include "bfm.sv"
`include "mon.sv"
`include "cov.sv"
`include "agent.sv"
`include "scb.sv"
`include "env.sv"
`include "assert.sv"
`include "tb.sv"

